`include "mux_5X1.v"
module tb();

	reg [4:0]i;
	reg [2:0]s;

	wire y;

	mux_5X1 dut(i,s,y);

	initial begin
		s=3'b000;i=5'b10000;#50;
		$display("s=%b i=%b y=%0d", s,i,y);

		s=3'b001;i=5'b01000;#50;
		$display("s=%b i=%b y=%0d", s,i,y);

		i=5'b11111;s=3'b010;#50;
		$display("s=%b i=%b y=%0d", s,i,y);

		s=3'b011;i=5'b00010;#50;
		$display("s=%b i=%b y=%0d", s,i,y);

		s=3'b100;i=5'b00001;#50;
		$display("s=%b i=%b y=%0d", s,i,y);


	end	

endmodule
